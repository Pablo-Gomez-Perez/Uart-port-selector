module main(input logic clk,
            input logic reset,
            input logic select,
            input logic Rx_ESP_Master,
            input logic Rx_Esp_Sim,
            input logic Rx_Pc_17,
            output logic Tx_Pc_18,
            output logic Tx_Esp_Master,
            output logic Tx_Esp_Sim,
            output logic Led_Selector);

    

endmodule